-- nios_cpu.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_cpu is
	port (
		clk_clk                                : in  std_logic                     := '0';             --                  clk.clk
		fpga_spi0_MISO                         : in  std_logic                     := '0';             --            fpga_spi0.MISO
		fpga_spi0_MOSI                         : out std_logic;                                        --                     .MOSI
		fpga_spi0_SCLK                         : out std_logic;                                        --                     .SCLK
		fpga_spi0_SS_n                         : out std_logic;                                        --                     .SS_n
		gpi0_export                            : in  std_logic_vector(7 downto 0)  := (others => '0'); --                 gpi0.export
		gpio0_export                           : out std_logic_vector(7 downto 0);                     --                gpio0.export
		pll_recfg_from_pll_0_reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => '0'); -- pll_recfg_from_pll_0.reconfig_from_pll
		pll_recfg_from_pll_1_reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => '0'); -- pll_recfg_from_pll_1.reconfig_from_pll
		pll_recfg_from_pll_2_reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => '0'); -- pll_recfg_from_pll_2.reconfig_from_pll
		pll_recfg_from_pll_3_reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => '0'); -- pll_recfg_from_pll_3.reconfig_from_pll
		pll_recfg_from_pll_4_reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => '0'); -- pll_recfg_from_pll_4.reconfig_from_pll
		pll_recfg_from_pll_5_reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => '0'); -- pll_recfg_from_pll_5.reconfig_from_pll
		pll_recfg_to_pll_0_reconfig_to_pll     : out std_logic_vector(63 downto 0);                    --   pll_recfg_to_pll_0.reconfig_to_pll
		pll_recfg_to_pll_1_reconfig_to_pll     : out std_logic_vector(63 downto 0);                    --   pll_recfg_to_pll_1.reconfig_to_pll
		pll_recfg_to_pll_2_reconfig_to_pll     : out std_logic_vector(63 downto 0);                    --   pll_recfg_to_pll_2.reconfig_to_pll
		pll_recfg_to_pll_3_reconfig_to_pll     : out std_logic_vector(63 downto 0);                    --   pll_recfg_to_pll_3.reconfig_to_pll
		pll_recfg_to_pll_4_reconfig_to_pll     : out std_logic_vector(63 downto 0);                    --   pll_recfg_to_pll_4.reconfig_to_pll
		pll_recfg_to_pll_5_reconfig_to_pll     : out std_logic_vector(63 downto 0);                    --   pll_recfg_to_pll_5.reconfig_to_pll
		pll_rst_export                         : out std_logic_vector(31 downto 0);                    --              pll_rst.export
		pllcfg_cmd_export                      : in  std_logic_vector(2 downto 0)  := (others => '0'); --           pllcfg_cmd.export
		pllcfg_spi_MISO                        : in  std_logic                     := '0';             --           pllcfg_spi.MISO
		pllcfg_spi_MOSI                        : out std_logic;                                        --                     .MOSI
		pllcfg_spi_SCLK                        : out std_logic;                                        --                     .SCLK
		pllcfg_spi_SS_n                        : out std_logic;                                        --                     .SS_n
		pllcfg_stat_export                     : out std_logic_vector(9 downto 0);                     --          pllcfg_stat.export
		reset_reset_n                          : out std_logic                                         --                reset.reset_n
	);
end entity nios_cpu;

architecture rtl of nios_cpu is
	component nios_cpu_PLLCFG_Command is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- export
		);
	end component nios_cpu_PLLCFG_Command;

	component nios_cpu_PLLCFG_SPI is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component nios_cpu_PLLCFG_SPI;

	component nios_cpu_PLLCFG_Status is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component nios_cpu_PLLCFG_Status;

	component nios_cpu_PLL_RST is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component nios_cpu_PLL_RST;

	component nios_cpu_fpga_spi0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component nios_cpu_fpga_spi0;

	component nios_cpu_gpi_0 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component nios_cpu_gpi_0;

	component nios_cpu_gpio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios_cpu_gpio_0;

	component nios_cpu_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_cpu_jtag_uart_0;

	component nios_cpu_nios2_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(15 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(15 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_cpu_nios2_cpu;

	component nios_cpu_oc_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios_cpu_oc_mem;

	component altera_pll_reconfig_top is
		generic (
			device_family       : string  := "";
			ENABLE_MIF          : boolean := false;
			MIF_FILE_NAME       : string  := "";
			ENABLE_BYTEENABLE   : boolean := false;
			BYTEENABLE_WIDTH    : integer := 4;
			RECONFIG_ADDR_WIDTH : integer := 6;
			RECONFIG_DATA_WIDTH : integer := 32;
			reconf_width        : integer := 64
		);
		port (
			mgmt_clk          : in  std_logic                     := 'X';             -- clk
			mgmt_reset        : in  std_logic                     := 'X';             -- reset
			mgmt_waitrequest  : out std_logic;                                        -- waitrequest
			mgmt_read         : in  std_logic                     := 'X';             -- read
			mgmt_write        : in  std_logic                     := 'X';             -- write
			mgmt_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			mgmt_address      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			mgmt_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reconfig_to_pll   : out std_logic_vector(63 downto 0);                    -- reconfig_to_pll
			reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => 'X'); -- reconfig_from_pll
			mgmt_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- byteenable
		);
	end component altera_pll_reconfig_top;

	component nios_cpu_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_cpu_sysid_qsys_0;

	component nios_cpu_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                : in  std_logic                     := 'X';             -- clk
			nios2_cpu_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			nios2_cpu_data_master_address                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios2_cpu_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			nios2_cpu_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_cpu_data_master_read                   : in  std_logic                     := 'X';             -- read
			nios2_cpu_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_cpu_data_master_write                  : in  std_logic                     := 'X';             -- write
			nios2_cpu_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_cpu_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			nios2_cpu_instruction_master_address         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios2_cpu_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			nios2_cpu_instruction_master_read            : in  std_logic                     := 'X';             -- read
			nios2_cpu_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			fpga_spi0_spi_control_port_address           : out std_logic_vector(2 downto 0);                     -- address
			fpga_spi0_spi_control_port_write             : out std_logic;                                        -- write
			fpga_spi0_spi_control_port_read              : out std_logic;                                        -- read
			fpga_spi0_spi_control_port_readdata          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			fpga_spi0_spi_control_port_writedata         : out std_logic_vector(15 downto 0);                    -- writedata
			fpga_spi0_spi_control_port_chipselect        : out std_logic;                                        -- chipselect
			gpi_0_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			gpi_0_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			gpio_0_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			gpio_0_s1_write                              : out std_logic;                                        -- write
			gpio_0_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			gpio_0_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			gpio_0_s1_chipselect                         : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address        : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write          : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read           : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest    : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect     : out std_logic;                                        -- chipselect
			nios2_cpu_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			nios2_cpu_debug_mem_slave_write              : out std_logic;                                        -- write
			nios2_cpu_debug_mem_slave_read               : out std_logic;                                        -- read
			nios2_cpu_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_cpu_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_cpu_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_cpu_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			nios2_cpu_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			oc_mem_s1_address                            : out std_logic_vector(11 downto 0);                    -- address
			oc_mem_s1_write                              : out std_logic;                                        -- write
			oc_mem_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			oc_mem_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			oc_mem_s1_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			oc_mem_s1_chipselect                         : out std_logic;                                        -- chipselect
			oc_mem_s1_clken                              : out std_logic;                                        -- clken
			pll_reconfig_0_mgmt_avalon_slave_address     : out std_logic_vector(5 downto 0);                     -- address
			pll_reconfig_0_mgmt_avalon_slave_write       : out std_logic;                                        -- write
			pll_reconfig_0_mgmt_avalon_slave_read        : out std_logic;                                        -- read
			pll_reconfig_0_mgmt_avalon_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_reconfig_0_mgmt_avalon_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			pll_reconfig_0_mgmt_avalon_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			pll_reconfig_1_mgmt_avalon_slave_address     : out std_logic_vector(5 downto 0);                     -- address
			pll_reconfig_1_mgmt_avalon_slave_write       : out std_logic;                                        -- write
			pll_reconfig_1_mgmt_avalon_slave_read        : out std_logic;                                        -- read
			pll_reconfig_1_mgmt_avalon_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_reconfig_1_mgmt_avalon_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			pll_reconfig_1_mgmt_avalon_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			pll_reconfig_2_mgmt_avalon_slave_address     : out std_logic_vector(5 downto 0);                     -- address
			pll_reconfig_2_mgmt_avalon_slave_write       : out std_logic;                                        -- write
			pll_reconfig_2_mgmt_avalon_slave_read        : out std_logic;                                        -- read
			pll_reconfig_2_mgmt_avalon_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_reconfig_2_mgmt_avalon_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			pll_reconfig_2_mgmt_avalon_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			pll_reconfig_3_mgmt_avalon_slave_address     : out std_logic_vector(5 downto 0);                     -- address
			pll_reconfig_3_mgmt_avalon_slave_write       : out std_logic;                                        -- write
			pll_reconfig_3_mgmt_avalon_slave_read        : out std_logic;                                        -- read
			pll_reconfig_3_mgmt_avalon_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_reconfig_3_mgmt_avalon_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			pll_reconfig_3_mgmt_avalon_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			pll_reconfig_4_mgmt_avalon_slave_address     : out std_logic_vector(5 downto 0);                     -- address
			pll_reconfig_4_mgmt_avalon_slave_write       : out std_logic;                                        -- write
			pll_reconfig_4_mgmt_avalon_slave_read        : out std_logic;                                        -- read
			pll_reconfig_4_mgmt_avalon_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_reconfig_4_mgmt_avalon_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			pll_reconfig_4_mgmt_avalon_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			pll_reconfig_5_mgmt_avalon_slave_address     : out std_logic_vector(5 downto 0);                     -- address
			pll_reconfig_5_mgmt_avalon_slave_write       : out std_logic;                                        -- write
			pll_reconfig_5_mgmt_avalon_slave_read        : out std_logic;                                        -- read
			pll_reconfig_5_mgmt_avalon_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_reconfig_5_mgmt_avalon_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			pll_reconfig_5_mgmt_avalon_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			PLL_RST_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			PLL_RST_s1_write                             : out std_logic;                                        -- write
			PLL_RST_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PLL_RST_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			PLL_RST_s1_chipselect                        : out std_logic;                                        -- chipselect
			PLLCFG_Command_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			PLLCFG_Command_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PLLCFG_SPI_spi_control_port_address          : out std_logic_vector(2 downto 0);                     -- address
			PLLCFG_SPI_spi_control_port_write            : out std_logic;                                        -- write
			PLLCFG_SPI_spi_control_port_read             : out std_logic;                                        -- read
			PLLCFG_SPI_spi_control_port_readdata         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			PLLCFG_SPI_spi_control_port_writedata        : out std_logic_vector(15 downto 0);                    -- writedata
			PLLCFG_SPI_spi_control_port_chipselect       : out std_logic;                                        -- chipselect
			PLLCFG_Status_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			PLLCFG_Status_s1_write                       : out std_logic;                                        -- write
			PLLCFG_Status_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PLLCFG_Status_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			PLLCFG_Status_s1_chipselect                  : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address           : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component nios_cpu_mm_interconnect_0;

	component nios_cpu_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_cpu_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_cpu_debug_reset_request_reset                             : std_logic;                     -- nios2_cpu:debug_reset_request -> [nios2_cpu_debug_reset_request_reset:in, rst_controller:reset_in0]
	signal nios2_cpu_data_master_readdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	signal nios2_cpu_data_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	signal nios2_cpu_data_master_debugaccess                               : std_logic;                     -- nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	signal nios2_cpu_data_master_address                                   : std_logic_vector(15 downto 0); -- nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	signal nios2_cpu_data_master_byteenable                                : std_logic_vector(3 downto 0);  -- nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	signal nios2_cpu_data_master_read                                      : std_logic;                     -- nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	signal nios2_cpu_data_master_write                                     : std_logic;                     -- nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	signal nios2_cpu_data_master_writedata                                 : std_logic_vector(31 downto 0); -- nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	signal nios2_cpu_instruction_master_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	signal nios2_cpu_instruction_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	signal nios2_cpu_instruction_master_address                            : std_logic_vector(15 downto 0); -- nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	signal nios2_cpu_instruction_master_read                               : std_logic;                     -- nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata            : std_logic_vector(31 downto 0); -- nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest         : std_logic;                     -- nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess         : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_address             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_read                : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_write               : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata     : std_logic_vector(31 downto 0); -- pll_reconfig_0:mgmt_readdata -> mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_readdata
	signal mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest  : std_logic;                     -- pll_reconfig_0:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_waitrequest
	signal mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address      : std_logic_vector(5 downto 0);  -- mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_address -> pll_reconfig_0:mgmt_address
	signal mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read         : std_logic;                     -- mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_read -> pll_reconfig_0:mgmt_read
	signal mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write        : std_logic;                     -- mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_write -> pll_reconfig_0:mgmt_write
	signal mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_writedata -> pll_reconfig_0:mgmt_writedata
	signal mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_readdata     : std_logic_vector(31 downto 0); -- pll_reconfig_5:mgmt_readdata -> mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_readdata
	signal mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_waitrequest  : std_logic;                     -- pll_reconfig_5:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_waitrequest
	signal mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_address      : std_logic_vector(5 downto 0);  -- mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_address -> pll_reconfig_5:mgmt_address
	signal mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_read         : std_logic;                     -- mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_read -> pll_reconfig_5:mgmt_read
	signal mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_write        : std_logic;                     -- mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_write -> pll_reconfig_5:mgmt_write
	signal mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_writedata -> pll_reconfig_5:mgmt_writedata
	signal mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_readdata     : std_logic_vector(31 downto 0); -- pll_reconfig_4:mgmt_readdata -> mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_readdata
	signal mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_waitrequest  : std_logic;                     -- pll_reconfig_4:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_waitrequest
	signal mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_address      : std_logic_vector(5 downto 0);  -- mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_address -> pll_reconfig_4:mgmt_address
	signal mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_read         : std_logic;                     -- mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_read -> pll_reconfig_4:mgmt_read
	signal mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_write        : std_logic;                     -- mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_write -> pll_reconfig_4:mgmt_write
	signal mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_writedata -> pll_reconfig_4:mgmt_writedata
	signal mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_readdata     : std_logic_vector(31 downto 0); -- pll_reconfig_3:mgmt_readdata -> mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_readdata
	signal mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_waitrequest  : std_logic;                     -- pll_reconfig_3:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_waitrequest
	signal mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_address      : std_logic_vector(5 downto 0);  -- mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_address -> pll_reconfig_3:mgmt_address
	signal mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_read         : std_logic;                     -- mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_read -> pll_reconfig_3:mgmt_read
	signal mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_write        : std_logic;                     -- mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_write -> pll_reconfig_3:mgmt_write
	signal mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_writedata -> pll_reconfig_3:mgmt_writedata
	signal mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_readdata     : std_logic_vector(31 downto 0); -- pll_reconfig_2:mgmt_readdata -> mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_readdata
	signal mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_waitrequest  : std_logic;                     -- pll_reconfig_2:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_waitrequest
	signal mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_address      : std_logic_vector(5 downto 0);  -- mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_address -> pll_reconfig_2:mgmt_address
	signal mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_read         : std_logic;                     -- mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_read -> pll_reconfig_2:mgmt_read
	signal mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_write        : std_logic;                     -- mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_write -> pll_reconfig_2:mgmt_write
	signal mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_writedata -> pll_reconfig_2:mgmt_writedata
	signal mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_readdata     : std_logic_vector(31 downto 0); -- pll_reconfig_1:mgmt_readdata -> mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_readdata
	signal mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_waitrequest  : std_logic;                     -- pll_reconfig_1:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_waitrequest
	signal mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_address      : std_logic_vector(5 downto 0);  -- mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_address -> pll_reconfig_1:mgmt_address
	signal mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_read         : std_logic;                     -- mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_read -> pll_reconfig_1:mgmt_read
	signal mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_write        : std_logic;                     -- mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_write -> pll_reconfig_1:mgmt_write
	signal mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_writedata -> pll_reconfig_1:mgmt_writedata
	signal mm_interconnect_0_oc_mem_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:oc_mem_s1_chipselect -> oc_mem:chipselect
	signal mm_interconnect_0_oc_mem_s1_readdata                            : std_logic_vector(31 downto 0); -- oc_mem:readdata -> mm_interconnect_0:oc_mem_s1_readdata
	signal mm_interconnect_0_oc_mem_s1_address                             : std_logic_vector(11 downto 0); -- mm_interconnect_0:oc_mem_s1_address -> oc_mem:address
	signal mm_interconnect_0_oc_mem_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:oc_mem_s1_byteenable -> oc_mem:byteenable
	signal mm_interconnect_0_oc_mem_s1_write                               : std_logic;                     -- mm_interconnect_0:oc_mem_s1_write -> oc_mem:write
	signal mm_interconnect_0_oc_mem_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:oc_mem_s1_writedata -> oc_mem:writedata
	signal mm_interconnect_0_oc_mem_s1_clken                               : std_logic;                     -- mm_interconnect_0:oc_mem_s1_clken -> oc_mem:clken
	signal mm_interconnect_0_gpio_0_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:gpio_0_s1_chipselect -> gpio_0:chipselect
	signal mm_interconnect_0_gpio_0_s1_readdata                            : std_logic_vector(31 downto 0); -- gpio_0:readdata -> mm_interconnect_0:gpio_0_s1_readdata
	signal mm_interconnect_0_gpio_0_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:gpio_0_s1_address -> gpio_0:address
	signal mm_interconnect_0_gpio_0_s1_write                               : std_logic;                     -- mm_interconnect_0:gpio_0_s1_write -> mm_interconnect_0_gpio_0_s1_write:in
	signal mm_interconnect_0_gpio_0_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:gpio_0_s1_writedata -> gpio_0:writedata
	signal mm_interconnect_0_gpi_0_s1_readdata                             : std_logic_vector(31 downto 0); -- gpi_0:readdata -> mm_interconnect_0:gpi_0_s1_readdata
	signal mm_interconnect_0_gpi_0_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:gpi_0_s1_address -> gpi_0:address
	signal mm_interconnect_0_pllcfg_command_s1_readdata                    : std_logic_vector(31 downto 0); -- PLLCFG_Command:readdata -> mm_interconnect_0:PLLCFG_Command_s1_readdata
	signal mm_interconnect_0_pllcfg_command_s1_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PLLCFG_Command_s1_address -> PLLCFG_Command:address
	signal mm_interconnect_0_pllcfg_status_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:PLLCFG_Status_s1_chipselect -> PLLCFG_Status:chipselect
	signal mm_interconnect_0_pllcfg_status_s1_readdata                     : std_logic_vector(31 downto 0); -- PLLCFG_Status:readdata -> mm_interconnect_0:PLLCFG_Status_s1_readdata
	signal mm_interconnect_0_pllcfg_status_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PLLCFG_Status_s1_address -> PLLCFG_Status:address
	signal mm_interconnect_0_pllcfg_status_s1_write                        : std_logic;                     -- mm_interconnect_0:PLLCFG_Status_s1_write -> mm_interconnect_0_pllcfg_status_s1_write:in
	signal mm_interconnect_0_pllcfg_status_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:PLLCFG_Status_s1_writedata -> PLLCFG_Status:writedata
	signal mm_interconnect_0_pll_rst_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:PLL_RST_s1_chipselect -> PLL_RST:chipselect
	signal mm_interconnect_0_pll_rst_s1_readdata                           : std_logic_vector(31 downto 0); -- PLL_RST:readdata -> mm_interconnect_0:PLL_RST_s1_readdata
	signal mm_interconnect_0_pll_rst_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PLL_RST_s1_address -> PLL_RST:address
	signal mm_interconnect_0_pll_rst_s1_write                              : std_logic;                     -- mm_interconnect_0:PLL_RST_s1_write -> mm_interconnect_0_pll_rst_s1_write:in
	signal mm_interconnect_0_pll_rst_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:PLL_RST_s1_writedata -> PLL_RST:writedata
	signal mm_interconnect_0_fpga_spi0_spi_control_port_chipselect         : std_logic;                     -- mm_interconnect_0:fpga_spi0_spi_control_port_chipselect -> fpga_spi0:spi_select
	signal mm_interconnect_0_fpga_spi0_spi_control_port_readdata           : std_logic_vector(15 downto 0); -- fpga_spi0:data_to_cpu -> mm_interconnect_0:fpga_spi0_spi_control_port_readdata
	signal mm_interconnect_0_fpga_spi0_spi_control_port_address            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:fpga_spi0_spi_control_port_address -> fpga_spi0:mem_addr
	signal mm_interconnect_0_fpga_spi0_spi_control_port_read               : std_logic;                     -- mm_interconnect_0:fpga_spi0_spi_control_port_read -> mm_interconnect_0_fpga_spi0_spi_control_port_read:in
	signal mm_interconnect_0_fpga_spi0_spi_control_port_write              : std_logic;                     -- mm_interconnect_0:fpga_spi0_spi_control_port_write -> mm_interconnect_0_fpga_spi0_spi_control_port_write:in
	signal mm_interconnect_0_fpga_spi0_spi_control_port_writedata          : std_logic_vector(15 downto 0); -- mm_interconnect_0:fpga_spi0_spi_control_port_writedata -> fpga_spi0:data_from_cpu
	signal mm_interconnect_0_pllcfg_spi_spi_control_port_chipselect        : std_logic;                     -- mm_interconnect_0:PLLCFG_SPI_spi_control_port_chipselect -> PLLCFG_SPI:spi_select
	signal mm_interconnect_0_pllcfg_spi_spi_control_port_readdata          : std_logic_vector(15 downto 0); -- PLLCFG_SPI:data_to_cpu -> mm_interconnect_0:PLLCFG_SPI_spi_control_port_readdata
	signal mm_interconnect_0_pllcfg_spi_spi_control_port_address           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:PLLCFG_SPI_spi_control_port_address -> PLLCFG_SPI:mem_addr
	signal mm_interconnect_0_pllcfg_spi_spi_control_port_read              : std_logic;                     -- mm_interconnect_0:PLLCFG_SPI_spi_control_port_read -> mm_interconnect_0_pllcfg_spi_spi_control_port_read:in
	signal mm_interconnect_0_pllcfg_spi_spi_control_port_write             : std_logic;                     -- mm_interconnect_0:PLLCFG_SPI_spi_control_port_write -> mm_interconnect_0_pllcfg_spi_spi_control_port_write:in
	signal mm_interconnect_0_pllcfg_spi_spi_control_port_writedata         : std_logic_vector(15 downto 0); -- mm_interconnect_0:PLLCFG_SPI_spi_control_port_writedata -> PLLCFG_SPI:data_from_cpu
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- fpga_spi0:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- PLLCFG_SPI:irq -> irq_mapper:receiver2_irq
	signal nios2_cpu_irq_irq                                               : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_cpu:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, oc_mem:reset, pll_reconfig_0:mgmt_reset, pll_reconfig_1:mgmt_reset, pll_reconfig_2:mgmt_reset, pll_reconfig_3:mgmt_reset, pll_reconfig_4:mgmt_reset, pll_reconfig_5:mgmt_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2_cpu:reset_req, oc_mem:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_gpio_0_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_gpio_0_s1_write:inv -> gpio_0:write_n
	signal mm_interconnect_0_pllcfg_status_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_pllcfg_status_s1_write:inv -> PLLCFG_Status:write_n
	signal mm_interconnect_0_pll_rst_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_pll_rst_s1_write:inv -> PLL_RST:write_n
	signal mm_interconnect_0_fpga_spi0_spi_control_port_read_ports_inv     : std_logic;                     -- mm_interconnect_0_fpga_spi0_spi_control_port_read:inv -> fpga_spi0:read_n
	signal mm_interconnect_0_fpga_spi0_spi_control_port_write_ports_inv    : std_logic;                     -- mm_interconnect_0_fpga_spi0_spi_control_port_write:inv -> fpga_spi0:write_n
	signal mm_interconnect_0_pllcfg_spi_spi_control_port_read_ports_inv    : std_logic;                     -- mm_interconnect_0_pllcfg_spi_spi_control_port_read:inv -> PLLCFG_SPI:read_n
	signal mm_interconnect_0_pllcfg_spi_spi_control_port_write_ports_inv   : std_logic;                     -- mm_interconnect_0_pllcfg_spi_spi_control_port_write:inv -> PLLCFG_SPI:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [PLLCFG_Command:reset_n, PLLCFG_SPI:reset_n, PLLCFG_Status:reset_n, PLL_RST:reset_n, fpga_spi0:reset_n, gpi_0:reset_n, gpio_0:reset_n, jtag_uart_0:rst_n, nios2_cpu:reset_n, sysid_qsys_0:reset_n]

begin

	pllcfg_command : component nios_cpu_PLLCFG_Command
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address  => mm_interconnect_0_pllcfg_command_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pllcfg_command_s1_readdata, --                    .readdata
			in_port  => pllcfg_cmd_export                             -- external_connection.export
		);

	pllcfg_spi : component nios_cpu_PLLCFG_SPI
		port map (
			clk           => clk_clk,                                                       --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                      --            reset.reset_n
			data_from_cpu => mm_interconnect_0_pllcfg_spi_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_pllcfg_spi_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_pllcfg_spi_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_pllcfg_spi_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_pllcfg_spi_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_pllcfg_spi_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver2_irq,                                      --              irq.irq
			MISO          => pllcfg_spi_MISO,                                               --         external.export
			MOSI          => pllcfg_spi_MOSI,                                               --                 .export
			SCLK          => pllcfg_spi_SCLK,                                               --                 .export
			SS_n          => pllcfg_spi_SS_n                                                --                 .export
		);

	pllcfg_status : component nios_cpu_PLLCFG_Status
		port map (
			clk        => clk_clk,                                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_pllcfg_status_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pllcfg_status_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pllcfg_status_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pllcfg_status_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pllcfg_status_s1_readdata,        --                    .readdata
			out_port   => pllcfg_stat_export                                  -- external_connection.export
		);

	pll_rst : component nios_cpu_PLL_RST
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pll_rst_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pll_rst_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pll_rst_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pll_rst_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pll_rst_s1_readdata,        --                    .readdata
			out_port   => pll_rst_export                                -- external_connection.export
		);

	fpga_spi0 : component nios_cpu_fpga_spi0
		port map (
			clk           => clk_clk,                                                      --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                     --            reset.reset_n
			data_from_cpu => mm_interconnect_0_fpga_spi0_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_fpga_spi0_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_fpga_spi0_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_fpga_spi0_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_fpga_spi0_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_fpga_spi0_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver1_irq,                                     --              irq.irq
			MISO          => fpga_spi0_MISO,                                               --         external.export
			MOSI          => fpga_spi0_MOSI,                                               --                 .export
			SCLK          => fpga_spi0_SCLK,                                               --                 .export
			SS_n          => fpga_spi0_SS_n                                                --                 .export
		);

	gpi_0 : component nios_cpu_gpi_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_gpi_0_s1_address,       --                  s1.address
			readdata => mm_interconnect_0_gpi_0_s1_readdata,      --                    .readdata
			in_port  => gpi0_export                               -- external_connection.export
		);

	gpio_0 : component nios_cpu_gpio_0
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_gpio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_gpio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_gpio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_gpio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_gpio_0_s1_readdata,        --                    .readdata
			out_port   => gpio0_export                                 -- external_connection.export
		);

	jtag_uart_0 : component nios_cpu_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	nios2_cpu : component nios_cpu_nios2_cpu
		port map (
			clk                                 => clk_clk,                                                 --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                      --                          .reset_req
			d_address                           => nios2_cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_cpu_data_master_read,                              --                          .read
			d_readdata                          => nios2_cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_cpu_data_master_write,                             --                          .write
			d_writedata                         => nios2_cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_cpu_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                     -- custom_instruction_master.readra
		);

	oc_mem : component nios_cpu_oc_mem
		port map (
			clk        => clk_clk,                                --   clk1.clk
			address    => mm_interconnect_0_oc_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_oc_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_oc_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_oc_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_oc_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_oc_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_oc_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,         -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req      --       .reset_req
		);

	pll_reconfig_0 : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64
		)
		port map (
			mgmt_clk          => clk_clk,                                                        --          mgmt_clk.clk
			mgmt_reset        => rst_controller_reset_out_reset,                                 --        mgmt_reset.reset
			mgmt_waitrequest  => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest, -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read,        --                  .read
			mgmt_write        => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write,       --                  .write
			mgmt_readdata     => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata,    --                  .readdata
			mgmt_address      => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address,     --                  .address
			mgmt_writedata    => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata,   --                  .writedata
			reconfig_to_pll   => pll_recfg_to_pll_0_reconfig_to_pll,                             --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => pll_recfg_from_pll_0_reconfig_from_pll,                         -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"                                                          --       (terminated)
		);

	pll_reconfig_1 : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64
		)
		port map (
			mgmt_clk          => clk_clk,                                                        --          mgmt_clk.clk
			mgmt_reset        => rst_controller_reset_out_reset,                                 --        mgmt_reset.reset
			mgmt_waitrequest  => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_waitrequest, -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_read,        --                  .read
			mgmt_write        => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_write,       --                  .write
			mgmt_readdata     => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_readdata,    --                  .readdata
			mgmt_address      => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_address,     --                  .address
			mgmt_writedata    => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_writedata,   --                  .writedata
			reconfig_to_pll   => pll_recfg_to_pll_1_reconfig_to_pll,                             --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => pll_recfg_from_pll_1_reconfig_from_pll,                         -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"                                                          --       (terminated)
		);

	pll_reconfig_2 : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64
		)
		port map (
			mgmt_clk          => clk_clk,                                                        --          mgmt_clk.clk
			mgmt_reset        => rst_controller_reset_out_reset,                                 --        mgmt_reset.reset
			mgmt_waitrequest  => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_waitrequest, -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_read,        --                  .read
			mgmt_write        => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_write,       --                  .write
			mgmt_readdata     => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_readdata,    --                  .readdata
			mgmt_address      => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_address,     --                  .address
			mgmt_writedata    => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_writedata,   --                  .writedata
			reconfig_to_pll   => pll_recfg_to_pll_2_reconfig_to_pll,                             --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => pll_recfg_from_pll_2_reconfig_from_pll,                         -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"                                                          --       (terminated)
		);

	pll_reconfig_3 : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64
		)
		port map (
			mgmt_clk          => clk_clk,                                                        --          mgmt_clk.clk
			mgmt_reset        => rst_controller_reset_out_reset,                                 --        mgmt_reset.reset
			mgmt_waitrequest  => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_waitrequest, -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_read,        --                  .read
			mgmt_write        => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_write,       --                  .write
			mgmt_readdata     => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_readdata,    --                  .readdata
			mgmt_address      => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_address,     --                  .address
			mgmt_writedata    => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_writedata,   --                  .writedata
			reconfig_to_pll   => pll_recfg_to_pll_3_reconfig_to_pll,                             --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => pll_recfg_from_pll_3_reconfig_from_pll,                         -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"                                                          --       (terminated)
		);

	pll_reconfig_4 : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64
		)
		port map (
			mgmt_clk          => clk_clk,                                                        --          mgmt_clk.clk
			mgmt_reset        => rst_controller_reset_out_reset,                                 --        mgmt_reset.reset
			mgmt_waitrequest  => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_waitrequest, -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_read,        --                  .read
			mgmt_write        => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_write,       --                  .write
			mgmt_readdata     => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_readdata,    --                  .readdata
			mgmt_address      => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_address,     --                  .address
			mgmt_writedata    => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_writedata,   --                  .writedata
			reconfig_to_pll   => pll_recfg_to_pll_4_reconfig_to_pll,                             --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => pll_recfg_from_pll_4_reconfig_from_pll,                         -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"                                                          --       (terminated)
		);

	pll_reconfig_5 : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64
		)
		port map (
			mgmt_clk          => clk_clk,                                                        --          mgmt_clk.clk
			mgmt_reset        => rst_controller_reset_out_reset,                                 --        mgmt_reset.reset
			mgmt_waitrequest  => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_waitrequest, -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_read,        --                  .read
			mgmt_write        => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_write,       --                  .write
			mgmt_readdata     => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_readdata,    --                  .readdata
			mgmt_address      => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_address,     --                  .address
			mgmt_writedata    => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_writedata,   --                  .writedata
			reconfig_to_pll   => pll_recfg_to_pll_5_reconfig_to_pll,                             --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => pll_recfg_from_pll_5_reconfig_from_pll,                         -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"                                                          --       (terminated)
		);

	sysid_qsys_0 : component nios_cpu_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component nios_cpu_mm_interconnect_0
		port map (
			clk_0_clk_clk                                => clk_clk,                                                        --                             clk_0_clk.clk
			nios2_cpu_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                                 -- nios2_cpu_reset_reset_bridge_in_reset.reset
			nios2_cpu_data_master_address                => nios2_cpu_data_master_address,                                  --                 nios2_cpu_data_master.address
			nios2_cpu_data_master_waitrequest            => nios2_cpu_data_master_waitrequest,                              --                                      .waitrequest
			nios2_cpu_data_master_byteenable             => nios2_cpu_data_master_byteenable,                               --                                      .byteenable
			nios2_cpu_data_master_read                   => nios2_cpu_data_master_read,                                     --                                      .read
			nios2_cpu_data_master_readdata               => nios2_cpu_data_master_readdata,                                 --                                      .readdata
			nios2_cpu_data_master_write                  => nios2_cpu_data_master_write,                                    --                                      .write
			nios2_cpu_data_master_writedata              => nios2_cpu_data_master_writedata,                                --                                      .writedata
			nios2_cpu_data_master_debugaccess            => nios2_cpu_data_master_debugaccess,                              --                                      .debugaccess
			nios2_cpu_instruction_master_address         => nios2_cpu_instruction_master_address,                           --          nios2_cpu_instruction_master.address
			nios2_cpu_instruction_master_waitrequest     => nios2_cpu_instruction_master_waitrequest,                       --                                      .waitrequest
			nios2_cpu_instruction_master_read            => nios2_cpu_instruction_master_read,                              --                                      .read
			nios2_cpu_instruction_master_readdata        => nios2_cpu_instruction_master_readdata,                          --                                      .readdata
			fpga_spi0_spi_control_port_address           => mm_interconnect_0_fpga_spi0_spi_control_port_address,           --            fpga_spi0_spi_control_port.address
			fpga_spi0_spi_control_port_write             => mm_interconnect_0_fpga_spi0_spi_control_port_write,             --                                      .write
			fpga_spi0_spi_control_port_read              => mm_interconnect_0_fpga_spi0_spi_control_port_read,              --                                      .read
			fpga_spi0_spi_control_port_readdata          => mm_interconnect_0_fpga_spi0_spi_control_port_readdata,          --                                      .readdata
			fpga_spi0_spi_control_port_writedata         => mm_interconnect_0_fpga_spi0_spi_control_port_writedata,         --                                      .writedata
			fpga_spi0_spi_control_port_chipselect        => mm_interconnect_0_fpga_spi0_spi_control_port_chipselect,        --                                      .chipselect
			gpi_0_s1_address                             => mm_interconnect_0_gpi_0_s1_address,                             --                              gpi_0_s1.address
			gpi_0_s1_readdata                            => mm_interconnect_0_gpi_0_s1_readdata,                            --                                      .readdata
			gpio_0_s1_address                            => mm_interconnect_0_gpio_0_s1_address,                            --                             gpio_0_s1.address
			gpio_0_s1_write                              => mm_interconnect_0_gpio_0_s1_write,                              --                                      .write
			gpio_0_s1_readdata                           => mm_interconnect_0_gpio_0_s1_readdata,                           --                                      .readdata
			gpio_0_s1_writedata                          => mm_interconnect_0_gpio_0_s1_writedata,                          --                                      .writedata
			gpio_0_s1_chipselect                         => mm_interconnect_0_gpio_0_s1_chipselect,                         --                                      .chipselect
			jtag_uart_0_avalon_jtag_slave_address        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,        --         jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,          --                                      .write
			jtag_uart_0_avalon_jtag_slave_read           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,           --                                      .read
			jtag_uart_0_avalon_jtag_slave_readdata       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,       --                                      .readdata
			jtag_uart_0_avalon_jtag_slave_writedata      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,      --                                      .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,    --                                      .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,     --                                      .chipselect
			nios2_cpu_debug_mem_slave_address            => mm_interconnect_0_nios2_cpu_debug_mem_slave_address,            --             nios2_cpu_debug_mem_slave.address
			nios2_cpu_debug_mem_slave_write              => mm_interconnect_0_nios2_cpu_debug_mem_slave_write,              --                                      .write
			nios2_cpu_debug_mem_slave_read               => mm_interconnect_0_nios2_cpu_debug_mem_slave_read,               --                                      .read
			nios2_cpu_debug_mem_slave_readdata           => mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata,           --                                      .readdata
			nios2_cpu_debug_mem_slave_writedata          => mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata,          --                                      .writedata
			nios2_cpu_debug_mem_slave_byteenable         => mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable,         --                                      .byteenable
			nios2_cpu_debug_mem_slave_waitrequest        => mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest,        --                                      .waitrequest
			nios2_cpu_debug_mem_slave_debugaccess        => mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess,        --                                      .debugaccess
			oc_mem_s1_address                            => mm_interconnect_0_oc_mem_s1_address,                            --                             oc_mem_s1.address
			oc_mem_s1_write                              => mm_interconnect_0_oc_mem_s1_write,                              --                                      .write
			oc_mem_s1_readdata                           => mm_interconnect_0_oc_mem_s1_readdata,                           --                                      .readdata
			oc_mem_s1_writedata                          => mm_interconnect_0_oc_mem_s1_writedata,                          --                                      .writedata
			oc_mem_s1_byteenable                         => mm_interconnect_0_oc_mem_s1_byteenable,                         --                                      .byteenable
			oc_mem_s1_chipselect                         => mm_interconnect_0_oc_mem_s1_chipselect,                         --                                      .chipselect
			oc_mem_s1_clken                              => mm_interconnect_0_oc_mem_s1_clken,                              --                                      .clken
			pll_reconfig_0_mgmt_avalon_slave_address     => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address,     --      pll_reconfig_0_mgmt_avalon_slave.address
			pll_reconfig_0_mgmt_avalon_slave_write       => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write,       --                                      .write
			pll_reconfig_0_mgmt_avalon_slave_read        => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read,        --                                      .read
			pll_reconfig_0_mgmt_avalon_slave_readdata    => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata,    --                                      .readdata
			pll_reconfig_0_mgmt_avalon_slave_writedata   => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata,   --                                      .writedata
			pll_reconfig_0_mgmt_avalon_slave_waitrequest => mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest, --                                      .waitrequest
			pll_reconfig_1_mgmt_avalon_slave_address     => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_address,     --      pll_reconfig_1_mgmt_avalon_slave.address
			pll_reconfig_1_mgmt_avalon_slave_write       => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_write,       --                                      .write
			pll_reconfig_1_mgmt_avalon_slave_read        => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_read,        --                                      .read
			pll_reconfig_1_mgmt_avalon_slave_readdata    => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_readdata,    --                                      .readdata
			pll_reconfig_1_mgmt_avalon_slave_writedata   => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_writedata,   --                                      .writedata
			pll_reconfig_1_mgmt_avalon_slave_waitrequest => mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_waitrequest, --                                      .waitrequest
			pll_reconfig_2_mgmt_avalon_slave_address     => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_address,     --      pll_reconfig_2_mgmt_avalon_slave.address
			pll_reconfig_2_mgmt_avalon_slave_write       => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_write,       --                                      .write
			pll_reconfig_2_mgmt_avalon_slave_read        => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_read,        --                                      .read
			pll_reconfig_2_mgmt_avalon_slave_readdata    => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_readdata,    --                                      .readdata
			pll_reconfig_2_mgmt_avalon_slave_writedata   => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_writedata,   --                                      .writedata
			pll_reconfig_2_mgmt_avalon_slave_waitrequest => mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_waitrequest, --                                      .waitrequest
			pll_reconfig_3_mgmt_avalon_slave_address     => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_address,     --      pll_reconfig_3_mgmt_avalon_slave.address
			pll_reconfig_3_mgmt_avalon_slave_write       => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_write,       --                                      .write
			pll_reconfig_3_mgmt_avalon_slave_read        => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_read,        --                                      .read
			pll_reconfig_3_mgmt_avalon_slave_readdata    => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_readdata,    --                                      .readdata
			pll_reconfig_3_mgmt_avalon_slave_writedata   => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_writedata,   --                                      .writedata
			pll_reconfig_3_mgmt_avalon_slave_waitrequest => mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_waitrequest, --                                      .waitrequest
			pll_reconfig_4_mgmt_avalon_slave_address     => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_address,     --      pll_reconfig_4_mgmt_avalon_slave.address
			pll_reconfig_4_mgmt_avalon_slave_write       => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_write,       --                                      .write
			pll_reconfig_4_mgmt_avalon_slave_read        => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_read,        --                                      .read
			pll_reconfig_4_mgmt_avalon_slave_readdata    => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_readdata,    --                                      .readdata
			pll_reconfig_4_mgmt_avalon_slave_writedata   => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_writedata,   --                                      .writedata
			pll_reconfig_4_mgmt_avalon_slave_waitrequest => mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_waitrequest, --                                      .waitrequest
			pll_reconfig_5_mgmt_avalon_slave_address     => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_address,     --      pll_reconfig_5_mgmt_avalon_slave.address
			pll_reconfig_5_mgmt_avalon_slave_write       => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_write,       --                                      .write
			pll_reconfig_5_mgmt_avalon_slave_read        => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_read,        --                                      .read
			pll_reconfig_5_mgmt_avalon_slave_readdata    => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_readdata,    --                                      .readdata
			pll_reconfig_5_mgmt_avalon_slave_writedata   => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_writedata,   --                                      .writedata
			pll_reconfig_5_mgmt_avalon_slave_waitrequest => mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_waitrequest, --                                      .waitrequest
			PLL_RST_s1_address                           => mm_interconnect_0_pll_rst_s1_address,                           --                            PLL_RST_s1.address
			PLL_RST_s1_write                             => mm_interconnect_0_pll_rst_s1_write,                             --                                      .write
			PLL_RST_s1_readdata                          => mm_interconnect_0_pll_rst_s1_readdata,                          --                                      .readdata
			PLL_RST_s1_writedata                         => mm_interconnect_0_pll_rst_s1_writedata,                         --                                      .writedata
			PLL_RST_s1_chipselect                        => mm_interconnect_0_pll_rst_s1_chipselect,                        --                                      .chipselect
			PLLCFG_Command_s1_address                    => mm_interconnect_0_pllcfg_command_s1_address,                    --                     PLLCFG_Command_s1.address
			PLLCFG_Command_s1_readdata                   => mm_interconnect_0_pllcfg_command_s1_readdata,                   --                                      .readdata
			PLLCFG_SPI_spi_control_port_address          => mm_interconnect_0_pllcfg_spi_spi_control_port_address,          --           PLLCFG_SPI_spi_control_port.address
			PLLCFG_SPI_spi_control_port_write            => mm_interconnect_0_pllcfg_spi_spi_control_port_write,            --                                      .write
			PLLCFG_SPI_spi_control_port_read             => mm_interconnect_0_pllcfg_spi_spi_control_port_read,             --                                      .read
			PLLCFG_SPI_spi_control_port_readdata         => mm_interconnect_0_pllcfg_spi_spi_control_port_readdata,         --                                      .readdata
			PLLCFG_SPI_spi_control_port_writedata        => mm_interconnect_0_pllcfg_spi_spi_control_port_writedata,        --                                      .writedata
			PLLCFG_SPI_spi_control_port_chipselect       => mm_interconnect_0_pllcfg_spi_spi_control_port_chipselect,       --                                      .chipselect
			PLLCFG_Status_s1_address                     => mm_interconnect_0_pllcfg_status_s1_address,                     --                      PLLCFG_Status_s1.address
			PLLCFG_Status_s1_write                       => mm_interconnect_0_pllcfg_status_s1_write,                       --                                      .write
			PLLCFG_Status_s1_readdata                    => mm_interconnect_0_pllcfg_status_s1_readdata,                    --                                      .readdata
			PLLCFG_Status_s1_writedata                   => mm_interconnect_0_pllcfg_status_s1_writedata,                   --                                      .writedata
			PLLCFG_Status_s1_chipselect                  => mm_interconnect_0_pllcfg_status_s1_chipselect,                  --                                      .chipselect
			sysid_qsys_0_control_slave_address           => mm_interconnect_0_sysid_qsys_0_control_slave_address,           --            sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata          => mm_interconnect_0_sysid_qsys_0_control_slave_readdata           --                                      .readdata
		);

	irq_mapper : component nios_cpu_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => nios2_cpu_irq_irq               --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_cpu_debug_reset_request_reset, -- reset_in0.reset
			clk            => clk_clk,                             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,  --          .reset_req
			reset_req_in0  => '0',                                 -- (terminated)
			reset_in1      => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	reset_reset_n <= not nios2_cpu_debug_reset_request_reset;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_gpio_0_s1_write_ports_inv <= not mm_interconnect_0_gpio_0_s1_write;

	mm_interconnect_0_pllcfg_status_s1_write_ports_inv <= not mm_interconnect_0_pllcfg_status_s1_write;

	mm_interconnect_0_pll_rst_s1_write_ports_inv <= not mm_interconnect_0_pll_rst_s1_write;

	mm_interconnect_0_fpga_spi0_spi_control_port_read_ports_inv <= not mm_interconnect_0_fpga_spi0_spi_control_port_read;

	mm_interconnect_0_fpga_spi0_spi_control_port_write_ports_inv <= not mm_interconnect_0_fpga_spi0_spi_control_port_write;

	mm_interconnect_0_pllcfg_spi_spi_control_port_read_ports_inv <= not mm_interconnect_0_pllcfg_spi_spi_control_port_read;

	mm_interconnect_0_pllcfg_spi_spi_control_port_write_ports_inv <= not mm_interconnect_0_pllcfg_spi_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_cpu
