LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY bypass IS

	GENERIC (N : NATURAL := 18);
	PORT (
		d : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
		q : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0));

END ENTITY bypass;

ARCHITECTURE beh OF bypass IS
BEGIN

	q <= d;

END ARCHITECTURE beh;